module Decoder(
    instr_op_i,
	RegWrite_o,
	ALU_op_o,
	ALUSrc_o,
	RegDst_o,
	Branch_o
	);

    //I/O ports
    input  [6-1:0] instr_op_i;

    output         RegWrite_o;
    output [3-1:0] ALU_op_o;
    output         ALUSrc_o;
    output         RegDst_o;
    output         Branch_o;

    //Internal Signals
    reg    [3-1:0] ALU_op_o;
    reg            ALUSrc_o;
    reg            RegWrite_o;
    reg            RegDst_o;
    reg            Branch_o;

    //Parameter


    //Main function
    always @ ( * ) begin
        if (instr_op_i == 6'b000000) begin      //r-type
            ALU_op_o  = 3'b010;
            ALUSrc_o  = 0;
            RegWrite_o= 1;
            RegDst_o  = 1;
            Branch_o  = 0;
        end
        else if (instr_op_i == 6'b110001) begin //lw
            ALU_op_o  = 3'b000;
            ALUSrc_o  = 1;
            RegWrite_o= 1;
            RegDst_o  = 0;
            Branch_o  = 0;
        end
        else if(instr_op_i == 6'b110101)begin  //sw
            ALU_op_o  = 3'b000;
            ALUSrc_o  = 1;
            RegWrite_o= 0;
            RegDst_o  = 1'bx;
            Branch_o  = 0;
        end
        else if(instr_op_i == 6'b001000)begin    //brench
            ALU_op_o   = 3'b001;
            ALUSrc_o   = 0;
            RegWrite_o = 0;
            RegDst_o   = 1'bx;
            Branch_o   = 1;
        end
        else begin
            ALU_op_o  = 3'bxxx;
            ALUSrc_o  = 1'bx;
            RegWrite_o= 1'bx;
            RegDst_o  = 1'bx;
            Branch_o  = 1'bx;
        end
    end
endmodule
